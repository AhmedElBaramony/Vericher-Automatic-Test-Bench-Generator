module mux_logical_tb;

  //INPUTS
    reg A;
   reg B;
   reg C;
   reg D;
   reg S;
   reg R;

  //OUTPUTS
    wire [2:0]O;

  //INISTANCE
  mux_logical T (.A (A),.B (B),.C (C),.D (D),.S (S),.R (R),.O (O));



  initial begin
    // Run the simulation for a specific time

    #10 A = 0;B = 0;C = 0;D = 0;S = 0;R = 0;
   #10 A = 0;B = 0;C = 0;D = 0;S = 0;R = 1;
   #10 A = 0;B = 0;C = 0;D = 0;S = 1;R = 0;
   #10 A = 0;B = 0;C = 0;D = 0;S = 1;R = 1;
   #10 A = 0;B = 0;C = 0;D = 1;S = 0;R = 0;
   #10 A = 0;B = 0;C = 0;D = 1;S = 0;R = 1;
   #10 A = 0;B = 0;C = 0;D = 1;S = 1;R = 0;
   #10 A = 0;B = 0;C = 0;D = 1;S = 1;R = 1;
   #10 A = 0;B = 0;C = 1;D = 0;S = 0;R = 0;
   #10 A = 0;B = 0;C = 1;D = 0;S = 0;R = 1;
   #10 A = 0;B = 0;C = 1;D = 0;S = 1;R = 0;
   #10 A = 0;B = 0;C = 1;D = 0;S = 1;R = 1;
   #10 A = 0;B = 0;C = 1;D = 1;S = 0;R = 0;
   #10 A = 0;B = 0;C = 1;D = 1;S = 0;R = 1;
   #10 A = 0;B = 0;C = 1;D = 1;S = 1;R = 0;
   #10 A = 0;B = 0;C = 1;D = 1;S = 1;R = 1;
   #10 A = 0;B = 1;C = 0;D = 0;S = 0;R = 0;
   #10 A = 0;B = 1;C = 0;D = 0;S = 0;R = 1;
   #10 A = 0;B = 1;C = 0;D = 0;S = 1;R = 0;
   #10 A = 0;B = 1;C = 0;D = 0;S = 1;R = 1;
   #10 A = 0;B = 1;C = 0;D = 1;S = 0;R = 0;
   #10 A = 0;B = 1;C = 0;D = 1;S = 0;R = 1;
   #10 A = 0;B = 1;C = 0;D = 1;S = 1;R = 0;
   #10 A = 0;B = 1;C = 0;D = 1;S = 1;R = 1;
   #10 A = 0;B = 1;C = 1;D = 0;S = 0;R = 0;
   #10 A = 0;B = 1;C = 1;D = 0;S = 0;R = 1;
   #10 A = 0;B = 1;C = 1;D = 0;S = 1;R = 0;
   #10 A = 0;B = 1;C = 1;D = 0;S = 1;R = 1;
   #10 A = 0;B = 1;C = 1;D = 1;S = 0;R = 0;
   #10 A = 0;B = 1;C = 1;D = 1;S = 0;R = 1;
   #10 A = 0;B = 1;C = 1;D = 1;S = 1;R = 0;
   #10 A = 0;B = 1;C = 1;D = 1;S = 1;R = 1;
   #10 A = 1;B = 0;C = 0;D = 0;S = 0;R = 0;
   #10 A = 1;B = 0;C = 0;D = 0;S = 0;R = 1;
   #10 A = 1;B = 0;C = 0;D = 0;S = 1;R = 0;
   #10 A = 1;B = 0;C = 0;D = 0;S = 1;R = 1;
   #10 A = 1;B = 0;C = 0;D = 1;S = 0;R = 0;
   #10 A = 1;B = 0;C = 0;D = 1;S = 0;R = 1;
   #10 A = 1;B = 0;C = 0;D = 1;S = 1;R = 0;
   #10 A = 1;B = 0;C = 0;D = 1;S = 1;R = 1;
   #10 A = 1;B = 0;C = 1;D = 0;S = 0;R = 0;
   #10 A = 1;B = 0;C = 1;D = 0;S = 0;R = 1;
   #10 A = 1;B = 0;C = 1;D = 0;S = 1;R = 0;
   #10 A = 1;B = 0;C = 1;D = 0;S = 1;R = 1;
   #10 A = 1;B = 0;C = 1;D = 1;S = 0;R = 0;
   #10 A = 1;B = 0;C = 1;D = 1;S = 0;R = 1;
   #10 A = 1;B = 0;C = 1;D = 1;S = 1;R = 0;
   #10 A = 1;B = 0;C = 1;D = 1;S = 1;R = 1;
   #10 A = 1;B = 1;C = 0;D = 0;S = 0;R = 0;
   #10 A = 1;B = 1;C = 0;D = 0;S = 0;R = 1;
   #10 A = 1;B = 1;C = 0;D = 0;S = 1;R = 0;
   #10 A = 1;B = 1;C = 0;D = 0;S = 1;R = 1;
   #10 A = 1;B = 1;C = 0;D = 1;S = 0;R = 0;
   #10 A = 1;B = 1;C = 0;D = 1;S = 0;R = 1;
   #10 A = 1;B = 1;C = 0;D = 1;S = 1;R = 0;
   #10 A = 1;B = 1;C = 0;D = 1;S = 1;R = 1;
   #10 A = 1;B = 1;C = 1;D = 0;S = 0;R = 0;
   #10 A = 1;B = 1;C = 1;D = 0;S = 0;R = 1;
   #10 A = 1;B = 1;C = 1;D = 0;S = 1;R = 0;
   #10 A = 1;B = 1;C = 1;D = 0;S = 1;R = 1;
   #10 A = 1;B = 1;C = 1;D = 1;S = 0;R = 0;
   #10 A = 1;B = 1;C = 1;D = 1;S = 0;R = 1;
   #10 A = 1;B = 1;C = 1;D = 1;S = 1;R = 0;
   #10 A = 1;B = 1;C = 1;D = 1;S = 1;R = 1;


    // End the simulation
    $stop;
  end

endmodule